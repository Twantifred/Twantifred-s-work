module bcd7seg(
	input       [3:0] data,           //输入:3位二进制
	output reg  [6:0] HEX0            //输出:3位二进制对应的数码管译码——>数字   
	);

always@ (*) begin
    case(data)
        4'b0000: HEX0=7'b0000_001;
        4'b0001: HEX0=7'b1001_111;
        4'b0010: HEX0=7'b0010_010;
        4'b0011: HEX0=7'b0000_110;

        4'b0100: HEX0=7'b1001_100;
        4'b0101: HEX0=7'b0100_100;
        4'b0110: HEX0=7'b0100_000;
        4'b0111: HEX0=7'b0001_111;

        4'b1000: HEX0=7'b0000_000;
        4'b1001: HEX0=7'b0000_100;
        4'b1010: HEX0=7'b0001_000;
        4'b1011: HEX0=7'b1100_000;
        
        4'b1100: HEX0=7'b0110_001;
        4'b1101: HEX0=7'b1000_010;
        4'b1110: HEX0=7'b0110_000;
        4'b1111: HEX0=7'b0111_000;
    endcase
end
endmodule
